* C:\Users\ASUS\OneDrive - American International University-Bangladesh\Desktop\Simulation\Schematic4.sch

* Schematics Version 9.1 - Web Update 1
* Sat Nov 26 22:49:33 2022



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic4.net"
.INC "Schematic4.als"


.probe


.END
