* C:\Users\ASUS\OneDrive - American International University-Bangladesh\Desktop\Simulation\Schematic7.sch

* Schematics Version 9.1 - Web Update 1
* Sat Nov 26 23:45:09 2022



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic7.net"
.INC "Schematic7.als"


.probe


.END
