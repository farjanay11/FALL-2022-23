* C:\Users\User\Desktop\IEC LAB PSPIECE Data & Schematics\Schematics\2.sch

* Schematics Version 9.1 - Web Update 1
* Sat Nov 26 23:25:29 2022



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "2.net"
.INC "2.als"


.probe


.END
