* C:\Users\User\Desktop\IEC LAB PSPIECE Data & Schematics\Schematics\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Sat Nov 26 23:06:37 2022



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
