* C:\Users\User\Desktop\IEC LAB PSPIECE Data & Schematics\Schematics\6.sch

* Schematics Version 9.1 - Web Update 1
* Sun Nov 27 00:41:07 2022



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "6.net"
.INC "6.als"


.probe


.END
