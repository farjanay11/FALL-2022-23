* C:\Users\User\Desktop\IEC LAB PSPIECE Data & Schematics\Schematics\Schematic0.1.sch

* Schematics Version 9.1 - Web Update 1
* Sat Nov 26 22:10:36 2022



** Analysis setup **
.tran 0ns 400ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic0.1.net"
.INC "Schematic0.1.als"


.probe


.END
