* C:\Users\ASUS\OneDrive - American International University-Bangladesh\Desktop\Iec Lab(\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Sat Nov 26 22:34:51 2022



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
