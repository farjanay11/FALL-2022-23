* C:\Users\ASUS\OneDrive - American International University-Bangladesh\Desktop\Simulation\Schematic3.sch

* Schematics Version 9.1 - Web Update 1
* Sat Nov 26 23:02:54 2022



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic3.net"
.INC "Schematic3.als"


.probe


.END
