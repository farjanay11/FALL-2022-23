* C:\Users\User\Desktop\IEC LAB PSPIECE Data & Schematics\Schematics\4.1.sch

* Schematics Version 9.1 - Web Update 1
* Sat Nov 26 23:52:29 2022



** Analysis setup **
.tran 0ns 200ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "4.1.net"
.INC "4.1.als"


.probe


.END
