* C:\Users\ASUS\OneDrive - American International University-Bangladesh\Desktop\Simulation\Schematic6.sch

* Schematics Version 9.1 - Web Update 1
* Sat Nov 26 23:28:18 2022



** Analysis setup **
.tran 0ns 50ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic6.net"
.INC "Schematic6.als"


.probe


.END
