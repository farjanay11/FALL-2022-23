* C:\Users\ASUS\OneDrive - American International University-Bangladesh\Desktop\Iec Lab(\Circuit8.sch

* Schematics Version 9.1 - Web Update 1
* Thu Nov 24 21:34:03 2022



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Circuit8.net"
.INC "Circuit8.als"


.probe


.END
