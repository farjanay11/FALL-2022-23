* C:\Users\User\Desktop\IEC LAB PSPIECE Data & Schematics\Schematics\7.sch

* Schematics Version 9.1 - Web Update 1
* Sun Nov 27 00:47:38 2022



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "7.net"
.INC "7.als"


.probe


.END
