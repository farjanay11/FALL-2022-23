* C:\Users\User\Desktop\IEC LAB PSPIECE Data & Schematics\Schematics\Schematic0.2.sch

* Schematics Version 9.1 - Web Update 1
* Sat Nov 26 22:52:00 2022



** Analysis setup **
.tran 0ns 40ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic0.2.net"
.INC "Schematic0.2.als"


.probe


.END
