* C:\Users\ASUS\OneDrive - American International University-Bangladesh\Desktop\IEC LAB PSPIECE Data & Schematics\Final Schematics\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Sun Dec 04 14:42:01 2022



** Analysis setup **
.tran 0ns 100ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
